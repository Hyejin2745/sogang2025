//------------------------------------------------------------------------------
// "amba_axi_lite_m6.v" generated for new I2C support, 2025-01-20
//------------------------------------------------------------------------------

module amba_axi_lite_m6
    #(parameter [31:0] P0_ADDR_START=32'h0_0000
     ,parameter [31:0] P1_ADDR_START=32'h1_0000
     ,parameter [31:0] P2_ADDR_START=32'h2_0000
     ,parameter [31:0] P3_ADDR_START=32'h3_0000
     ,parameter [31:0] P4_ADDR_START=32'h4_0000
     ,parameter [31:0] P5_ADDR_START=32'h5_0000
     ,parameter [31:0] P0_SIZE=32'h1_0000
     ,parameter [31:0] P1_SIZE=32'h1_0000
     ,parameter [31:0] P2_SIZE=32'h1_0000
     ,parameter [31:0] P3_SIZE=32'h1_0000
     ,parameter [31:0] P4_SIZE=32'h1_0000
     ,parameter [31:0] P5_SIZE=32'h1_0000)
(
    input  wire        axi_lite_aresetn,
    input  wire        axi_lite_aclk   ,

    input  wire [31:0] s_axi_lite_awaddr ,
    input  wire        s_axi_lite_awvalid,
    output wire        s_axi_lite_awready,
    input  wire [31:0] s_axi_lite_wdata  ,
    input  wire        s_axi_lite_wvalid ,
    output wire        s_axi_lite_wready ,
    output wire [ 1:0] s_axi_lite_bresp  ,
    output wire        s_axi_lite_bvalid ,
    input  wire        s_axi_lite_bready ,
    input  wire [31:0] s_axi_lite_araddr ,
    input  wire        s_axi_lite_arvalid,
    output wire        s_axi_lite_arready,
    output wire [31:0] s_axi_lite_rdata  ,
    output wire [ 1:0] s_axi_lite_rresp  ,
    output wire        s_axi_lite_rvalid ,
    input  wire        s_axi_lite_rready ,
    output reg  [31:0] m0_axi_lite_awaddr ,
    output reg         m0_axi_lite_awvalid,
    input  wire        m0_axi_lite_awready,
    output reg  [31:0] m0_axi_lite_wdata  ,
    output reg         m0_axi_lite_wvalid ,
    input  wire        m0_axi_lite_wready ,
    input  wire [ 1:0] m0_axi_lite_bresp  ,
    input  wire        m0_axi_lite_bvalid ,
    output reg         m0_axi_lite_bready ,
    output reg  [31:0] m0_axi_lite_araddr ,
    output reg         m0_axi_lite_arvalid,
    input  wire        m0_axi_lite_arready,
    input  wire [31:0] m0_axi_lite_rdata  ,
    input  wire [ 1:0] m0_axi_lite_rresp  ,
    input  wire        m0_axi_lite_rvalid ,
    output reg         m0_axi_lite_rready ,
    output reg  [31:0] m1_axi_lite_awaddr ,
    output reg         m1_axi_lite_awvalid,
    input  wire        m1_axi_lite_awready,
    output reg  [31:0] m1_axi_lite_wdata  ,
    output reg         m1_axi_lite_wvalid ,
    input  wire        m1_axi_lite_wready ,
    input  wire [ 1:0] m1_axi_lite_bresp  ,
    input  wire        m1_axi_lite_bvalid ,
    output reg         m1_axi_lite_bready ,
    output reg  [31:0] m1_axi_lite_araddr ,
    output reg         m1_axi_lite_arvalid,
    input  wire        m1_axi_lite_arready,
    input  wire [31:0] m1_axi_lite_rdata  ,
    input  wire [ 1:0] m1_axi_lite_rresp  ,
    input  wire        m1_axi_lite_rvalid ,
    output reg         m1_axi_lite_rready ,
    output reg  [31:0] m2_axi_lite_awaddr ,
    output reg         m2_axi_lite_awvalid,
    input  wire        m2_axi_lite_awready,
    output reg  [31:0] m2_axi_lite_wdata  ,
    output reg         m2_axi_lite_wvalid ,
    input  wire        m2_axi_lite_wready ,
    input  wire [ 1:0] m2_axi_lite_bresp  ,
    input  wire        m2_axi_lite_bvalid ,
    output reg         m2_axi_lite_bready ,
    output reg  [31:0] m2_axi_lite_araddr ,
    output reg         m2_axi_lite_arvalid,
    input  wire        m2_axi_lite_arready,
    input  wire [31:0] m2_axi_lite_rdata  ,
    input  wire [ 1:0] m2_axi_lite_rresp  ,
    input  wire        m2_axi_lite_rvalid ,
    output reg         m2_axi_lite_rready ,
    output reg  [31:0] m3_axi_lite_awaddr ,
    output reg         m3_axi_lite_awvalid,
    input  wire        m3_axi_lite_awready,
    output reg  [31:0] m3_axi_lite_wdata  ,
    output reg         m3_axi_lite_wvalid ,
    input  wire        m3_axi_lite_wready ,
    input  wire [ 1:0] m3_axi_lite_bresp  ,
    input  wire        m3_axi_lite_bvalid ,
    output reg         m3_axi_lite_bready ,
    output reg  [31:0] m3_axi_lite_araddr ,
    output reg         m3_axi_lite_arvalid,
    input  wire        m3_axi_lite_arready,
    input  wire [31:0] m3_axi_lite_rdata  ,
    input  wire [ 1:0] m3_axi_lite_rresp  ,
    input  wire        m3_axi_lite_rvalid ,
    output reg         m3_axi_lite_rready ,
    output reg  [31:0] m4_axi_lite_awaddr ,
    output reg         m4_axi_lite_awvalid,
    input  wire        m4_axi_lite_awready,
    output reg  [31:0] m4_axi_lite_wdata  ,
    output reg         m4_axi_lite_wvalid ,
    input  wire        m4_axi_lite_wready ,
    input  wire [ 1:0] m4_axi_lite_bresp  ,
    input  wire        m4_axi_lite_bvalid ,
    output reg         m4_axi_lite_bready ,
    output reg  [31:0] m4_axi_lite_araddr ,
    output reg         m4_axi_lite_arvalid,
    input  wire        m4_axi_lite_arready,
    input  wire [31:0] m4_axi_lite_rdata  ,
    input  wire [ 1:0] m4_axi_lite_rresp  ,
    input  wire        m4_axi_lite_rvalid ,
    output reg         m4_axi_lite_rready ,
    output reg  [31:0] m5_axi_lite_awaddr ,
    output reg         m5_axi_lite_awvalid,
    input  wire        m5_axi_lite_awready,
    output reg  [31:0] m5_axi_lite_wdata  ,
    output reg         m5_axi_lite_wvalid ,
    input  wire        m5_axi_lite_wready ,
    input  wire [ 1:0] m5_axi_lite_bresp  ,
    input  wire        m5_axi_lite_bvalid ,
    output reg         m5_axi_lite_bready ,
    output reg  [31:0] m5_axi_lite_araddr ,
    output reg         m5_axi_lite_arvalid,
    input  wire        m5_axi_lite_arready,
    input  wire [31:0] m5_axi_lite_rdata  ,
    input  wire [ 1:0] m5_axi_lite_rresp  ,
    input  wire        m5_axi_lite_rvalid ,
    output reg         m5_axi_lite_rready  
);
    localparam [6*32-1:0] P_ADDR_START={P5_ADDR_START,P4_ADDR_START,P3_ADDR_START,P2_ADDR_START,P1_ADDR_START,P0_ADDR_START};
    localparam [6*32-1:0] P_SIZE={P5_SIZE,P4_SIZE,P3_SIZE,P2_SIZE,P1_SIZE,P0_SIZE};
    wire [6*32-1:0] m_axi_lite_awaddr ;
    wire [6-1:0]    m_axi_lite_awvalid;
    reg  [6-1:0]    m_axi_lite_awready;
    wire [6*32-1:0] m_axi_lite_wdata  ;
    wire [6-1:0]    m_axi_lite_wvalid ;
    reg  [6-1:0]    m_axi_lite_wready ;
    reg  [6*2-1:0]  m_axi_lite_bresp  ;
    reg  [6-1:0]    m_axi_lite_bvalid ;
    wire [6-1:0]    m_axi_lite_bready ;
    wire [6*32-1:0] m_axi_lite_araddr ;
    wire [6-1:0]    m_axi_lite_arvalid;
    reg  [6-1:0]    m_axi_lite_arready;
    reg  [6*32-1:0] m_axi_lite_rdata  ;
    reg  [6*2-1:0]  m_axi_lite_rresp  ;
    reg  [6-1:0]    m_axi_lite_rvalid ;
    wire [6-1:0]    m_axi_lite_rready ;
    always @ ( * ) begin
        m0_axi_lite_awaddr                 = m_axi_lite_awaddr       [32*0+:32];
        m0_axi_lite_awvalid                = m_axi_lite_awvalid      [0];
        m_axi_lite_awready      [0]        = m0_axi_lite_awready;
        m0_axi_lite_wdata                  = m_axi_lite_wdata        [32*0+:32];
        m0_axi_lite_wvalid                 = m_axi_lite_wvalid       [0];
        m_axi_lite_wready       [0]        = m0_axi_lite_wready ;
        m_axi_lite_bresp        [2*0+:2]   = m0_axi_lite_bresp  ;
        m_axi_lite_bvalid       [0]        = m0_axi_lite_bvalid ;
        m0_axi_lite_bready                 = m_axi_lite_bready       [0];
        m0_axi_lite_araddr                 = m_axi_lite_araddr       [32*0+:32];
        m0_axi_lite_arvalid                = m_axi_lite_arvalid      [0];
        m_axi_lite_arready      [0]        = m0_axi_lite_arready;
        m_axi_lite_rdata        [32*0+:32] = m0_axi_lite_rdata  ;
        m_axi_lite_rresp        [2*0+:2]   = m0_axi_lite_rresp  ;
        m_axi_lite_rvalid       [0]        = m0_axi_lite_rvalid ;
        m0_axi_lite_rready                 = m_axi_lite_rready       [0];
        m1_axi_lite_awaddr                 = m_axi_lite_awaddr       [32*1+:32];
        m1_axi_lite_awvalid                = m_axi_lite_awvalid      [1];
        m_axi_lite_awready      [1]        = m1_axi_lite_awready;
        m1_axi_lite_wdata                  = m_axi_lite_wdata        [32*1+:32];
        m1_axi_lite_wvalid                 = m_axi_lite_wvalid       [1];
        m_axi_lite_wready       [1]        = m1_axi_lite_wready ;
        m_axi_lite_bresp        [2*1+:2]   = m1_axi_lite_bresp  ;
        m_axi_lite_bvalid       [1]        = m1_axi_lite_bvalid ;
        m1_axi_lite_bready                 = m_axi_lite_bready       [1];
        m1_axi_lite_araddr                 = m_axi_lite_araddr       [32*1+:32];
        m1_axi_lite_arvalid                = m_axi_lite_arvalid      [1];
        m_axi_lite_arready      [1]        = m1_axi_lite_arready;
        m_axi_lite_rdata        [32*1+:32] = m1_axi_lite_rdata  ;
        m_axi_lite_rresp        [2*1+:2]   = m1_axi_lite_rresp  ;
        m_axi_lite_rvalid       [1]        = m1_axi_lite_rvalid ;
        m1_axi_lite_rready                 = m_axi_lite_rready       [1];
        m2_axi_lite_awaddr                 = m_axi_lite_awaddr       [32*2+:32];
        m2_axi_lite_awvalid                = m_axi_lite_awvalid      [2];
        m_axi_lite_awready      [2]        = m2_axi_lite_awready;
        m2_axi_lite_wdata                  = m_axi_lite_wdata        [32*2+:32];
        m2_axi_lite_wvalid                 = m_axi_lite_wvalid       [2];
        m_axi_lite_wready       [2]        = m2_axi_lite_wready ;
        m_axi_lite_bresp        [2*2+:2]   = m2_axi_lite_bresp  ;
        m_axi_lite_bvalid       [2]        = m2_axi_lite_bvalid ;
        m2_axi_lite_bready                 = m_axi_lite_bready       [2];
        m2_axi_lite_araddr                 = m_axi_lite_araddr       [32*2+:32];
        m2_axi_lite_arvalid                = m_axi_lite_arvalid      [2];
        m_axi_lite_arready      [2]        = m2_axi_lite_arready;
        m_axi_lite_rdata        [32*2+:32] = m2_axi_lite_rdata  ;
        m_axi_lite_rresp        [2*2+:2]   = m2_axi_lite_rresp  ;
        m_axi_lite_rvalid       [2]        = m2_axi_lite_rvalid ;
        m2_axi_lite_rready                 = m_axi_lite_rready       [2];
        m3_axi_lite_awaddr                 = m_axi_lite_awaddr       [32*3+:32];
        m3_axi_lite_awvalid                = m_axi_lite_awvalid      [3];
        m_axi_lite_awready      [3]        = m3_axi_lite_awready;
        m3_axi_lite_wdata                  = m_axi_lite_wdata        [32*3+:32];
        m3_axi_lite_wvalid                 = m_axi_lite_wvalid       [3];
        m_axi_lite_wready       [3]        = m3_axi_lite_wready ;
        m_axi_lite_bresp        [2*3+:2]   = m3_axi_lite_bresp  ;
        m_axi_lite_bvalid       [3]        = m3_axi_lite_bvalid ;
        m3_axi_lite_bready                 = m_axi_lite_bready       [3];
        m3_axi_lite_araddr                 = m_axi_lite_araddr       [32*3+:32];
        m3_axi_lite_arvalid                = m_axi_lite_arvalid      [3];
        m_axi_lite_arready      [3]        = m3_axi_lite_arready;
        m_axi_lite_rdata        [32*3+:32] = m3_axi_lite_rdata  ;
        m_axi_lite_rresp        [2*3+:2]   = m3_axi_lite_rresp  ;
        m_axi_lite_rvalid       [3]        = m3_axi_lite_rvalid ;
        m3_axi_lite_rready                 = m_axi_lite_rready       [3];
        m4_axi_lite_awaddr                 = m_axi_lite_awaddr       [32*4+:32];
        m4_axi_lite_awvalid                = m_axi_lite_awvalid      [4];
        m_axi_lite_awready      [4]        = m4_axi_lite_awready;
        m4_axi_lite_wdata                  = m_axi_lite_wdata        [32*4+:32];
        m4_axi_lite_wvalid                 = m_axi_lite_wvalid       [4];
        m_axi_lite_wready       [4]        = m4_axi_lite_wready ;
        m_axi_lite_bresp        [2*4+:2]   = m4_axi_lite_bresp  ;
        m_axi_lite_bvalid       [4]        = m4_axi_lite_bvalid ;
        m4_axi_lite_bready                 = m_axi_lite_bready       [4];
        m4_axi_lite_araddr                 = m_axi_lite_araddr       [32*4+:32];
        m4_axi_lite_arvalid                = m_axi_lite_arvalid      [4];
        m_axi_lite_arready      [4]        = m4_axi_lite_arready;
        m_axi_lite_rdata        [32*4+:32] = m4_axi_lite_rdata  ;
        m_axi_lite_rresp        [2*4+:2]   = m4_axi_lite_rresp  ;
        m_axi_lite_rvalid       [4]        = m4_axi_lite_rvalid ;
        m4_axi_lite_rready                 = m_axi_lite_rready       [4];
        m5_axi_lite_awaddr                 = m_axi_lite_awaddr       [32*5+:32];
        m5_axi_lite_awvalid                = m_axi_lite_awvalid      [5];
        m_axi_lite_awready      [5]        = m5_axi_lite_awready;
        m5_axi_lite_wdata                  = m_axi_lite_wdata        [32*5+:32];
        m5_axi_lite_wvalid                 = m_axi_lite_wvalid       [5];
        m_axi_lite_wready       [5]        = m5_axi_lite_wready ;
        m_axi_lite_bresp        [2*5+:2]   = m5_axi_lite_bresp  ;
        m_axi_lite_bvalid       [5]        = m5_axi_lite_bvalid ;
        m5_axi_lite_bready                 = m_axi_lite_bready       [5];
        m5_axi_lite_araddr                 = m_axi_lite_araddr       [32*5+:32];
        m5_axi_lite_arvalid                = m_axi_lite_arvalid      [5];
        m_axi_lite_arready      [5]        = m5_axi_lite_arready;
        m_axi_lite_rdata        [32*5+:32] = m5_axi_lite_rdata  ;
        m_axi_lite_rresp        [2*5+:2]   = m5_axi_lite_rresp  ;
        m_axi_lite_rvalid       [5]        = m5_axi_lite_rvalid ;
        m5_axi_lite_rready                 = m_axi_lite_rready       [5];
    end
    amba_axi_lite_m6_core #(.P_NUM_MST   (6  )
                        ,.P_ADDR_START(P_ADDR_START)
                        ,.P_SIZE      (P_SIZE      ))
    u_amba_axi_lite_m6_core (
          .axi_lite_aresetn   ( axi_lite_aresetn   )
        , .axi_lite_aclk      ( axi_lite_aclk      )
        , .s_axi_lite_awaddr  ( s_axi_lite_awaddr  )
        , .s_axi_lite_awvalid ( s_axi_lite_awvalid )
        , .s_axi_lite_awready ( s_axi_lite_awready )
        , .s_axi_lite_wdata   ( s_axi_lite_wdata   )
        , .s_axi_lite_wvalid  ( s_axi_lite_wvalid  )
        , .s_axi_lite_wready  ( s_axi_lite_wready  )
        , .s_axi_lite_bresp   ( s_axi_lite_bresp   )
        , .s_axi_lite_bvalid  ( s_axi_lite_bvalid  )
        , .s_axi_lite_bready  ( s_axi_lite_bready  )
        , .s_axi_lite_araddr  ( s_axi_lite_araddr  )
        , .s_axi_lite_arvalid ( s_axi_lite_arvalid )
        , .s_axi_lite_arready ( s_axi_lite_arready )
        , .s_axi_lite_rdata   ( s_axi_lite_rdata   )
        , .s_axi_lite_rresp   ( s_axi_lite_rresp   )
        , .s_axi_lite_rvalid  ( s_axi_lite_rvalid  )
        , .s_axi_lite_rready  ( s_axi_lite_rready  )
        , .m_axi_lite_awaddr  ( m_axi_lite_awaddr  )
        , .m_axi_lite_awvalid ( m_axi_lite_awvalid )
        , .m_axi_lite_awready ( m_axi_lite_awready )
        , .m_axi_lite_wdata   ( m_axi_lite_wdata   )
        , .m_axi_lite_wvalid  ( m_axi_lite_wvalid  )
        , .m_axi_lite_wready  ( m_axi_lite_wready  )
        , .m_axi_lite_bresp   ( m_axi_lite_bresp   )
        , .m_axi_lite_bvalid  ( m_axi_lite_bvalid  )
        , .m_axi_lite_bready  ( m_axi_lite_bready  )
        , .m_axi_lite_araddr  ( m_axi_lite_araddr  )
        , .m_axi_lite_arvalid ( m_axi_lite_arvalid )
        , .m_axi_lite_arready ( m_axi_lite_arready )
        , .m_axi_lite_rdata   ( m_axi_lite_rdata   )
        , .m_axi_lite_rresp   ( m_axi_lite_rresp   )
        , .m_axi_lite_rvalid  ( m_axi_lite_rvalid  )
        , .m_axi_lite_rready  ( m_axi_lite_rready  )
    );
endmodule
`ifndef amba_axi_lite_m6_CORE_V
`define amba_axi_lite_m6_CORE_V
//------------------------------------------------------------------------------
//  Copyright (c) 2023-2024 by Ando Ki.
//  All right reserved.
//
//  All rights are reserved by Ando Ki.
//------------------------------------------------------------------------------

module amba_axi_lite_m6_core
     #(parameter integer P_NUM_MST=6
      ,parameter [P_NUM_MST*32-1:0] P_ADDR_START={P_NUM_MST{32'h0000_0000}}
      ,parameter [P_NUM_MST*32-1:0] P_SIZE ={P_NUM_MST{32'h0001_0000}})
(
    input  wire       axi_lite_aresetn,
    input  wire       axi_lite_aclk   ,

    input  wire [31:0] s_axi_lite_awaddr ,
    input  wire        s_axi_lite_awvalid,
    output reg         s_axi_lite_awready,
    input  wire [31:0] s_axi_lite_wdata  ,
    input  wire        s_axi_lite_wvalid ,
    output reg         s_axi_lite_wready ,
    output reg  [ 1:0] s_axi_lite_bresp  ,
    output reg         s_axi_lite_bvalid ,
    input  wire        s_axi_lite_bready ,
    input  wire [31:0] s_axi_lite_araddr ,
    input  wire        s_axi_lite_arvalid,
    output reg         s_axi_lite_arready,
    output reg  [31:0] s_axi_lite_rdata  ,
    output reg  [ 1:0] s_axi_lite_rresp  ,
    output reg         s_axi_lite_rvalid ,
    input  wire        s_axi_lite_rready ,

    output reg  [P_NUM_MST*32-1:0]  m_axi_lite_awaddr ,
    output reg  [P_NUM_MST-1:0]     m_axi_lite_awvalid,
    input  wire [P_NUM_MST-1:0]     m_axi_lite_awready,
    output reg  [P_NUM_MST*32-1:0]  m_axi_lite_wdata  ,
    output reg  [P_NUM_MST-1:0]     m_axi_lite_wvalid ,
    input  wire [P_NUM_MST-1:0]     m_axi_lite_wready ,
    input  wire [P_NUM_MST*2-1:0]   m_axi_lite_bresp  ,
    input  wire [P_NUM_MST-1:0]     m_axi_lite_bvalid ,
    output reg  [P_NUM_MST-1:0]     m_axi_lite_bready ,
    output reg  [P_NUM_MST*32-1:0]  m_axi_lite_araddr ,
    output reg  [P_NUM_MST-1:0]     m_axi_lite_arvalid,
    input  wire [P_NUM_MST-1:0]     m_axi_lite_arready,
    input  wire [P_NUM_MST*32-1:0]  m_axi_lite_rdata  ,
    input  wire [P_NUM_MST*2-1:0]   m_axi_lite_rresp  ,
    input  wire [P_NUM_MST-1:0]     m_axi_lite_rvalid ,
    output reg  [P_NUM_MST-1:0]     m_axi_lite_rready
);
    //--------------------------------------------------------------------------
    reg  [31:0]  axil_awaddr ;
    reg          axil_awvalid;
    reg          axil_awready;
    reg  [31:0]  axil_wdata  ;
    reg          axil_wvalid ;
    reg          axil_wready ;
    reg  [ 1:0]  axil_bresp  ;
    reg          axil_bvalid ;
    reg          axil_bready ;
    //--------------------------------------------------------------------------
    localparam P_BITS=(P_NUM_MST);
    reg  [P_BITS-1:0] sel_write='h0;
    wire [P_BITS:0]   decoder_write=decoder(s_axi_lite_awaddr);
    //--------------------------------------------------------------------------
    localparam STW_ADDR ='h0
             , STW_DATA ='h1
             , STW_RESP ='h2
             , STW_ERROR='h3
             , STW_END  ='h4;
    reg [3:0] stateW=STW_ADDR;
    //--------------------------------------------------------------------------
    always @ (posedge axi_lite_aclk or negedge axi_lite_aresetn) begin
    if (axi_lite_aresetn==1'b0) begin
        axil_awaddr  <=  'h0;
        axil_awvalid <= 1'b0;
        axil_wdata   <=  'h0;
        axil_wvalid  <= 1'b0;
        axil_bready  <= 1'b0;
        s_axi_lite_awready <= 1'b0;
        s_axi_lite_wready  <= 1'b0;
        s_axi_lite_bresp   <=  'h0;
        s_axi_lite_bvalid  <= 1'b0;
        sel_write          <=  'h0;
        stateW             <= STW_ADDR;
    end else begin
    case (stateW)
    STW_ADDR: begin
        s_axi_lite_awready <= 1'b1;
        if (s_axi_lite_awvalid&s_axi_lite_awready) begin
            if (decoder_write[P_BITS]) begin
              axil_awaddr  <= 32'h0;
              axil_awvalid <= 1'b0;
              s_axi_lite_awready <= 1'b0;
              s_axi_lite_wready  <= 1'b1;
              sel_write    <= decoder_write[P_BITS-1:0];
              stateW       <= STW_ERROR;
            end else begin
              s_axi_lite_awready <= 1'b0;
              axil_awaddr  <= s_axi_lite_awaddr;
              axil_awvalid <= 1'b1;
              sel_write    <= decoder_write[P_BITS-1:0];
              stateW       <= STW_DATA;
            end
        end
        end // STW_ADDR
    STW_DATA: begin
        if (axil_awready) begin
            axil_awvalid      <= 1'b0;
            s_axi_lite_wready <= 1'b1;
        end
        if (s_axi_lite_wvalid&s_axi_lite_wready) begin
            s_axi_lite_wready <= 1'b0;
            axil_wdata  <= s_axi_lite_wdata;
            axil_wvalid <= 1'b1;
            stateW      <= STW_RESP;
        end
        end // STW_DATA
    STW_RESP: begin
        if (axil_wready) begin
            axil_wvalid <= 1'b0;
            axil_bready <= 1'b1;
        end
        if (axil_bvalid&axil_bready) begin
            axil_bready       <= 1'b0;
            s_axi_lite_bresp  <= axil_bresp;
            s_axi_lite_bvalid <= 1'b1;
            stateW            <= STW_END;
        end
        end // STW_RESP
    STW_ERROR: begin
        if (s_axi_lite_wvalid&s_axi_lite_wready) begin
            s_axi_lite_wready <= 1'b0;
            s_axi_lite_bresp  <=  2'b11; // decoder error
            s_axi_lite_bvalid <=  1'b1;
            stateW            <= STW_END;
        end
        end // STW_ERROR
    STW_END: begin
        if (s_axi_lite_bvalid&s_axi_lite_bready) begin
            s_axi_lite_bvalid  <= 1'b0;
            s_axi_lite_awready <= 1'b1;
            stateW             <= STW_ADDR;
        end
        end // STW_END
    default: begin
        axil_awaddr  <=  'h0;
        axil_awvalid <= 1'b0;
        axil_wdata   <=  'h0;
        axil_wvalid  <= 1'b0;
        axil_bready  <= 1'b0;
        s_axi_lite_bresp  <=  'h0;
        s_axi_lite_bvalid <= 1'b0;
        stateW            <= STW_ADDR;
             end
    endcase
    end // if
    end // always
    //--------------------------------------------------------------------------
    always @ ( * ) begin
        m_axi_lite_awaddr  = 32'h0;
        m_axi_lite_awvalid =  1'b0;
        m_axi_lite_wdata   = 32'h0;
        m_axi_lite_wvalid  =  1'b0;
        m_axi_lite_bready  =  1'b0;

        m_axi_lite_awaddr [sel_write*32+:32] = axil_awaddr ;
        m_axi_lite_awvalid[sel_write]        = axil_awvalid;
        m_axi_lite_wdata  [sel_write*32+:32] = axil_wdata  ;
        m_axi_lite_wvalid [sel_write]        = axil_wvalid ;
        m_axi_lite_bready [sel_write]        = axil_bready ;

        axil_awready = m_axi_lite_awready[sel_write];
        axil_wready  = m_axi_lite_wready [sel_write];
        axil_bresp   = m_axi_lite_bresp  [sel_write*2+:2];
        axil_bvalid  = m_axi_lite_bvalid [sel_write];
    end
    //--------------------------------------------------------------------------
    // synthesis translate_off
    reg  [8*20-1:0] stateW_ascii="ADDR";
    always @ (stateW) begin
    case (stateW)
     STW_ADDR : stateW_ascii="ADDR ";
     STW_DATA : stateW_ascii="DATA ";
     STW_RESP : stateW_ascii="DATA ";
     STW_ERROR: stateW_ascii="ERROR";
     STW_END  : stateW_ascii="END  ";
    default   : stateW_ascii="Unknown";
    endcase
    end // always
    // synthesis translate_on
    //--------------------------------------------------------------------------
    reg  [31:0]  axil_araddr ;
    reg          axil_arvalid;
    reg          axil_arready;
    reg  [31:0]  axil_rdata  ;
    reg  [ 1:0]  axil_rresp  ;
    reg          axil_rvalid ;
    reg          axil_rready ;
    //--------------------------------------------------------------------------
    reg  [P_BITS-1:0] sel_read='h0;
    wire [P_BITS  :0] decoder_read=decoder(s_axi_lite_araddr);
    //--------------------------------------------------------------------------
    localparam STR_ADDR ='h0
             , STR_DATA ='h1
             , STR_ERROR='h2
             , STR_END  ='h3;
    reg [1:0] stateR=STR_ADDR;
    //--------------------------------------------------------------------------
    always @ (posedge axi_lite_aclk or negedge axi_lite_aresetn) begin
    if (axi_lite_aresetn==1'b0) begin
        axil_araddr  <=  'h0;
        axil_arvalid <= 1'b0;
        axil_rready  <= 1'b0;
        s_axi_lite_arready <= 1'b0;
        s_axi_lite_rdata   <=  'h0;
        s_axi_lite_rresp   <= 2'b00;
        s_axi_lite_rvalid  <= 1'b0;
        stateR             <= STR_ADDR;
    end else begin
    case (stateR)
    STR_ADDR: begin
        s_axi_lite_arready <= 1'b1;
        if (s_axi_lite_arvalid&s_axi_lite_arready) begin
            if (decoder_read[P_BITS]) begin
                axil_araddr  <= 32'h0;
                axil_arvalid <=  1'b0;
                sel_read <= decoder_read[P_BITS-1:0];
                s_axi_lite_arready <= 1'b0;
                stateR       <= STR_ERROR;
            end else begin
                axil_araddr  <= s_axi_lite_araddr;
                axil_arvalid <= 1'b1;
                sel_read <= decoder_read[P_BITS-1:0];
                s_axi_lite_arready <= 1'b0;
                stateR   <= STR_DATA;
            end
        end
        end // STR_ADDR
    STR_DATA: begin
        if (axil_arready) begin
            axil_arvalid <= 1'b0;
            axil_rready  <= 1'b1;
        end
        if (axil_rvalid&axil_rready) begin
            axil_rready       <= 1'b0;
            s_axi_lite_rdata  <= axil_rdata;
            s_axi_lite_rresp  <= 2'b00;
            s_axi_lite_rvalid <= 1'b1;
            stateR            <= STR_END;
        end
        end // STR_DATA
    STR_ERROR: begin
        axil_rready       <=  1'b0;
        s_axi_lite_rdata  <= 32'h0;
        s_axi_lite_rresp  <=  2'b11; // decoder error
        s_axi_lite_rvalid <=  1'b1;
        stateR            <= STR_END;
        end // STR_ERROR
    STR_END: begin
        if (s_axi_lite_rvalid&s_axi_lite_rready) begin
            s_axi_lite_rvalid <= 1'b0;
            stateR            <= STR_ADDR;
        end
        end // STR_END
    default: begin
        axil_araddr  <=  'h0;
        axil_arvalid <= 1'b0;
        s_axi_lite_arready <= 1'b1;
        s_axi_lite_rresp   <=  'h0;
        s_axi_lite_rvalid  <= 1'b0;
        stateR             <= STR_ADDR;
             end
    endcase
    end // if
    end // always
    //--------------------------------------------------------------------------
    always @ ( * ) begin
        m_axi_lite_araddr  = 32'h0;
        m_axi_lite_arvalid =  1'b0;
        m_axi_lite_rready  =  1'b0;

        m_axi_lite_araddr [sel_read*32+:32] = axil_araddr ;
        m_axi_lite_arvalid[sel_read] = axil_arvalid;
        m_axi_lite_rready [sel_read] = axil_rready ;

        axil_arready = m_axi_lite_arready[sel_read];
        axil_rdata   = m_axi_lite_rdata  [sel_read*32+:32];
        axil_rresp   = m_axi_lite_rresp  [sel_read*2+:2];
        axil_rvalid  = m_axi_lite_rvalid [sel_read];
    end
    //--------------------------------------------------------------------------
    // synthesis translate_off
    reg  [8*20-1:0] stateR_ascii="ADDR";
    always @ (stateR) begin
    case (stateR)
     STR_ADDR : stateR_ascii="ADDR ";
     STR_DATA : stateR_ascii="DATA ";
     STR_ERROR: stateR_ascii="ERROR";
     STR_END  : stateR_ascii="END  ";
    default   : stateR_ascii="Unknown";
    endcase
    end // always
    // synthesis translate_on
    //--------------------------------------------------------------------------
    function [P_BITS:0] decoder;
        input [31:0] addr;
        reg [P_NUM_MST-1:0] sel;
        integer idx, idy;
    begin
        decoder = {1'b1, {P_BITS{1'b0}}}; // default
        for (idx=P_NUM_MST-1; idx>=0; idx=idx-1) begin
             if ((addr>=P_ADDR_START[idx*32+:32])&&
                 (addr<(P_ADDR_START[idx*32+:32]+P_SIZE[idx*32+:32])))
                  decoder = {1'b0,idx[P_BITS-1:0]};
        end
    end
    endfunction
    //--------------------------------------------------------------------------
    // synthesis translate_off
    integer idx, idy;
    reg [31:0] startX, startY;
    reg [31:0] endX, endY;
    initial begin
        for (idx=0; idx<P_NUM_MST; idx=idx+1) begin
             if (P_SIZE[idx*32+:32]=='h0) begin
                 $display("%m ERROR %0d address space zero.", idx);
             end
             startX = P_ADDR_START[idx*32+:32];
             endX = P_ADDR_START[idx*32+:32]+P_SIZE[idx*32+:32]-1;
        for (idy=idx+1; idy<P_NUM_MST; idy=idy+1) begin
             startY = P_ADDR_START[idy*32+:32];
             endY = P_ADDR_START[idy*32+:32]+P_SIZE[idy*32+:32]-1;
             if (((startX>=startY)&&(startX<=endY))||
                 ((endX  >=startY)&&(endX  <=endY))||
                 ((startY>=startX)&&(startY<=endX))||
                 ((endY  >=startX)&&(endY  <=endX))) begin
                 $display("%m ERROR address overlapped %0d:%0d.", idx, idy);
                 $display("\t[%0d]0x%08X-0x%08X [%0d]0x%08X-0x%08X", idx, startX, endX, idy, startY, endY);
             end
        end
        end
    end
    // synthesis translate_on
    //--------------------------------------------------------------------------
endmodule

//------------------------------------------------------------------------------
// Revision History
//
// 2025.01.20: Updated by Ando Ki (andoki@gmail.com) for new I2C support
//------------------------------------------------------------------------------
`endif // amba_axi_lite_m6_CORE_V

